module ysyx_24120013_top(
    input clk,
    input rst
);

endmodule