`timescale 1ns / 1ps
module top(
    input clk,
    input rst
);

endmodule