module ysyx_24120013_PC (
    input clk,
    input rst,
    input clear_en,
    output reg[31:0] pc
);

always @(posedge clk) begin
    ;
end

endmodule