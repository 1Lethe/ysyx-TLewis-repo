module ysyx_24120013_RegisterFile #(ADDR_WIDTH = 5, DATA_WIDTH = 32) (
        input clk,
        input rst,
        input [DATA_WIDTH-1:0] wdata,
        input [ADDR_WIDTH-1:0] waddr,
        input wen,
        input [ADDR_WIDTH-1:0] raddr1,
        input [ADDR_WIDTH-1:0] raddr2,
        output wire [DATA_WIDTH-1:0] rdata1,
        output wire [DATA_WIDTH-1:0] rdata2,

        output wire [DATA_WIDTH-1:0] rf_dis [2**ADDR_WIDTH-1:0],
        output wire [DATA_WIDTH-1:0] trap_flag
    );

    reg [DATA_WIDTH-1:0] rf [2**ADDR_WIDTH-1:0];

    always @(posedge clk) begin
        if(wen) begin
            rf[waddr] <= wdata;
        end
        rf[0] <= {DATA_WIDTH{1'b0}};
    end

    assign rdata1 = rf[raddr1];
    assign rdata2 = rf[raddr2];

    assign rf_dis = rf;
    assign trap_flag = rf[10];

endmodule
