module ysyx_24120013_top(
    input clk,
    input rst,
    input [31:0] pmem
);

endmodule